* File: DFFPOSX1.pex.netlist
* Created: Wed Jan  2 18:36:24 2008
* Program "Calibre xRC"
* Version "v2007.2_34.24"
* 
.subckt dff D Q clk vdd gnd
* 
MM21 Q a_66_6# gnd gnd nch L=5e-08 W=5e-07
MM19 a_76_6# a_2_6# a_66_6# gnd nch L=5e-08 W=2.5e-07
MM20 gnd Q a_76_6# gnd nch L=5e-08 W=2.5e-07
MM18 a_66_6# clk a_61_6# gnd nch L=5e-08 W=2.5e-07
MM17 a_61_6# a_34_4# gnd gnd nch L=5e-08 W=2.5e-07
MM10 gnd clk a_2_6# gnd nch L=5e-08 W=5e-07
MM16 a_34_4# a_22_6# gnd gnd nch L=5e-08 W=2.5e-07
MM15 gnd a_34_4# a_31_6# gnd nch L=5e-08 W=2.5e-07
MM14 a_31_6# clk a_22_6# gnd nch L=5e-08 W=2.5e-07
MM13 a_22_6# a_2_6# a_17_6# gnd nch L=5e-08 W=2.5e-07
MM12 a_17_6# D gnd gnd nch L=5e-08 W=2.5e-07
MM11 Q a_66_6# vdd vdd pch L=5e-08 W=1e-06
MM9 vdd Q a_76_84# vdd pch L=5e-08 W=2.5e-07
MM8 a_76_84# clk a_66_6# vdd pch L=5e-08 W=2.5e-07
MM7 a_66_6# a_2_6# a_61_74# vdd pch L=5e-08 W=5e-07
MM6 a_61_74# a_34_4# vdd vdd pch L=5e-08 W=5e-07
MM0 vdd clk a_2_6# vdd pch L=5e-08 W=1e-06
MM5 a_34_4# a_22_6# vdd vdd pch L=5e-08 W=5e-07
MM4 vdd a_34_4# a_31_74# vdd pch L=5e-08 W=5e-07
MM3 a_31_74# a_2_6# a_22_6# vdd pch L=5e-08 W=5e-07
MM2 a_22_6# clk a_17_74# vdd pch L=5e-08 W=5e-07
MM1 a_17_74# D vdd vdd pch L=5e-08 W=5e-07
* c_9 a_66_6# 0 0.271997f
* c_20 clk 0 0.350944f
* c_27 Q 0 0.202617f
* c_32 a_76_84# 0 0.0210573f
* c_38 a_76_6# 0 0.0204911f
* c_45 a_34_4# 0 0.172306f
* c_55 a_2_6# 0 0.283119f
* c_59 a_22_6# 0 0.157312f
* c_64 D 0 0.0816386f
* c_73 gnd 0 0.254131f
* c_81 vdd 0 0.23624f
*
*.include "dff.pex.netlist.dff.pxi"
*
.ends
*
*

.subckt replica_os_gc rbl wbl rwl wwl vdd
xi4 rbl vdd rwl osfet W=120e-9
xi3 wbl wwl vdd osfet W=70e-9
.ends replica_os_gc
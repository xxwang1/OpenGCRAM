
.SUBCKT tri_gate in out en en_bar vdd gnd
M_1 net_2 in_inv gnd gnd nch_mac W=180.000000n L=50.000000n
M_2 out en net_2 gnd nch_mac W=180.000000n L=50.000000n
M_3 net_3 in_inv vdd vdd pch_mac W=360.000000n L=50.000000n
M_4 out en_bar net_3 vdd pch_mac W=360.000000n L=50.000000n
M_5 in_inv in vdd vdd pch_mac W=180.000000n L=50.000000n
M_6 in_inv in gnd gnd nch_mac W=90.000000n L=50.000000n
.ENDS


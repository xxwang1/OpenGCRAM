
.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pch w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nch w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pch w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nch w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pch w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pch w=360.000000n l=50.000000n
mout0N bl en int2 gnd nch w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nch w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pch w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pch w=360.000000n l=50.000000n
mout1N br en int4 gnd nch w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nch w=180.000000n l=50.000000n
.ENDS write_driver


.subckt dummy_os_gc rbl wbl rwl wwl
xi4 rbl_noconn sn rwl osfet W=120e-9
xi3 wbl_noconn wwl sn osfet W=70e-9
.ends dummy_os_gc
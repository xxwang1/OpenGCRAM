.subckt os_gc rbl wbl rwl wwl
xi4 rbl sn rwl osfet W=120e-9
xi3 wbl wwl sn osfet W=70e-9
.ends os_gc